library IEEE;
use ieee.numeric_bit.all;

entity log_fd is

end log_fd;

architecture arch of log_fd is
end architecture;
