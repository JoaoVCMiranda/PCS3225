library IEEE;

