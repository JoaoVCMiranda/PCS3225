library IEEE;
use ieee.numeric_bit.all;

entity log_uc is

end log_uc;

architecture arch of log_uc is
end architecture;
